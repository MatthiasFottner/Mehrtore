* C:\Users\David\Documents\Studium\GitHub\UE Elektrische Netzwerke und Mehrtore\Mehrtore\UE_3\PSpice\Schalterposition a\Schalterposition a.sch

* Schematics Version 9.1 - Web Update 1
* Tue Nov 10 17:02:41 2020



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schalterposition a.net"
.INC "Schalterposition a.als"


.probe


.END
