** Profile: "SCHEMATIC1-uebung1"  [ C:\Users\matth\OneDrive - Technische Universit�t Graz\Dokumente\Studium\Graz\Semester_3\Elektrische_Netzwerke_und_Mehrtore\UE\UE_1\PSpice\erweitertes_KSV\simulation-SCHEMATIC1-uebung1.sim ] 

** Creating circuit file "simulation-SCHEMATIC1-uebung1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of pspiceev.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.PROBE 
.INC "simulation-SCHEMATIC1.net" 

.INC "simulation-SCHEMATIC1.als"


.END
