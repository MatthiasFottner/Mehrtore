* C:\Users\matth\OneDrive - Technische Universit�t Graz\Dokumente\Studium\Graz\Semester_3\Elektrische_Netzwerke_und_Mehrtore\UE_git\UE_2\PSpice\GR04_UE_02_whole_circuit_original.sch

* Schematics Version 9.1 - Web Update 1
* Mon Nov 02 22:48:21 2020



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "GR04_UE_02_whole_circuit_original.net"
.INC "GR04_UE_02_whole_circuit_original.als"


.probe


.END
