* C:\Users\David\Documents\Studium\GitHub\UE Elektrische Netzwerke und Mehrtore\Mehrtore\UE_3\PSpice\Testschematic.sch

* Schematics Version 9.1 - Web Update 1
* Sun Nov 08 15:39:14 2020



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Testschematic.net"
.INC "Testschematic.als"


.probe


.END
